1|1|x|s|0|assets\|realms_vernon|
1|1|x|s|0|assets\|realms_natalis|
1|1|x|s|0|assets\|realms_esterad|
1|0|1|s|0|assets\|realms_redania|
1|0|1|s|0|assets\|realms_redania_1|
1|0|1|s|0|assets\|realms_poor_infantry|
1|0|1|s|0|assets\|realms_poor_infantry|
1|0|1|s|0|assets\|realms_poor_infantry|
1|0|2|s|0|assets\|realms_yarpen|
1|0|4|s|0|assets\|realms_blue_stripes|
1|0|4|s|0|assets\|realms_blue_stripes|
1|0|4|s|0|assets\|realms_blue_stripes|
1|0|4|s|0|assets\|realms_dijkstra|
1|0|5|s|0|assets\|realms_ves|
1|0|5|s|0|assets\|realms_stennis|
1|0|5|s|0|assets\|realms_siegfried|
1|1|x|b|0|assets\|realms_philippa|
1|0|4|b|0|assets\|realms_sabrina|
1|0|4|b|0|assets\|realms_sheldon|
1|0|5|b|0|assets\|realms_keira|
1|0|5|b|0|assets\|realms_crinfrid|
1|0|5|b|0|assets\|realms_crinfrid|
1|0|5|b|0|assets\|realms_crinfrid|
1|0|5|b|0|assets\|realms_sheala|
1|0|6|b|0|assets\|realms_dethmold|
1|0|1|a|0|assets\|realms_kaedwen_siege|
1|0|1|a|0|assets\|realms_kaedwen_siege_1|
1|0|1|a|0|assets\|realms_kaedwen_siege_2|
1|0|1|a|0|assets\|realms_thaler|
1|0|5|a|0|assets\|realms_banner_nurse|
1|0|6|a|0|assets\|realms_ballista|
1|0|6|a|0|assets\|realms_trebuchet|
1|0|6|a|0|assets\|realms_siege_tower|
1|0|8|a|0|assets\|realms_catapult_1|
1|0|8|a|0|assets\|realms_catapult_1|
2|1|x|s|0|assets\|nilfgaard_letho|
2|1|x|s|0|assets\|nilfgaard_menno|
2|0|2|s|0|assets\|nilfgaard_vreemde|
2|0|2|s|0|assets\|nilfgaard_nauzicaa_2|
2|0|2|s|0|assets\|nilfgaard_nauzicaa_2|
2|0|2|s|0|assets\|nilfgaard_nauzicaa_2|
2|0|3|s|0|assets\|nilfgaard_imperal_brigade|
2|0|3|s|0|assets\|nilfgaard_imperal_brigade|
2|0|3|s|0|assets\|nilfgaard_imperal_brigade|
2|0|3|s|0|assets\|nilfgaard_morteisen|
2|0|4|s|0|assets\|nilfgaard_vattier|
2|0|4|s|0|assets\|nilfgaard_rainfarn|
2|0|5|s|0|assets\|nilfgaard_young_emissary|
2|0|5|s|0|assets\|nilfgaard_young_emissary_1|
2|0|6|s|0|assets\|nilfgaard_cahir|
2|0|7|s|0|assets\|nilfgaard_shilard|
2|0|9|s|0|assets\|nilfgaard_stefan|
2|1|x|b|0|assets\|nilfgaard_tibor|
2|0|1|b|0|assets\|nilfgaard_archer_support|
2|0|1|b|0|assets\|nilfgaard_archer_support_1|
2|0|1|b|0|assets\|nilfgaard_archer_support_1|
2|0|2|b|0|assets\|nilfgaard_albrich|
2|0|2|b|0|assets\|nilfgaard_sweers|
2|0|3|b|0|assets\|nilfgaard_puttkammer|
2|0|4|b|0|assets\|nilfgaard_vanhemar|
2|0|4|b|0|assets\|nilfgaard_cynthia|
2|0|5|b|0|assets\|nilfgaard_renuald|
2|0|6|b|0|assets\|nilfgaard_assire|
2|0|6|b|0|assets\|nilfgaard_fringilla|
2|0|x|b|0|assets\|nilfgaard_black_archer|
2|1|x|a|0|assets\|nilfgaard_moorvran|
2|0|0|a|0|assets\|nilfgaard_siege_support|
2|0|3|a|0|assets\|nilfgaard_rotten|
2|0|5|a|0|assets\|nilfgaard_zerri|
2|0|x|a|0|assets\|nilfgaard_heavy_zerri|
0|1|0|s|0|assets\|neutral_mysterious_elf|
0|1|7|s|0|assets\|neutral_triss|
0|1|l|s|0|assets\|neutral_geralt|
0|1|l|s|0|assets\|neutral_ciri|
0|0|2|s|0|assets\|neutral_dandelion|
0|0|5|s|0|assets\|neutral_zoltan|
0|0|5|s|0|assets\|neutral_emiel|
0|0|6|s|0|assets\|neutral_vesemir|
0|0|7|s|0|assets\|neutral_villen|
0|1|7|b|0|assets\|neutral_yennefer|