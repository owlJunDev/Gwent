Player|0|0|